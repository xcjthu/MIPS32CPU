// Module:  mem_wb
// File:    mem_wb.v
// Description: MEM/WB�׶εļĴ���
// Revision: 1.0
//////////////////////////////////////////////////////////////////////

`include "defines.v"

module mem_wb(

	input wire clk,
	input wire rst,
	

	//���Էô�׶ε���Ϣ	
	input wire[`RegAddrBus]       mem_wd,
	input wire                    mem_wreg,
	input wire[`RegBus]           mem_wdata,

	//�͵���д�׶ε���Ϣ
	output reg[`RegAddrBus]      wb_wd,
	output reg                   wb_wreg,
    output reg[`RegBus]          wb_wdata	       
	
);


	always @ (posedge clk) begin
		if(rst == `RstEnable) begin
			wb_wd <= `NOPRegAddr;
			wb_wreg <= `WriteDisable;
		  wb_wdata <= `ZeroWord;	
		end else begin
			wb_wd <= mem_wd;
			wb_wreg <= mem_wreg;
			wb_wdata <= mem_wdata;
		end    //if
	end      //always
			

endmodule